module div(rs1_reg,rs2_reg);
endmodule
